
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create a pulse for A 
*Va A VGND pulse(0 1.8 1n 10p 10p 1n 2n)
Va0 A0 VGND pulse(0   1.8 1000p 10p 10p 1000p 2000p)
Va1 A1 VGND pulse(1.8 0   1000p 10p 10p 1000p 2000p)
Vs  S  VGND pulse(0   1.8 500p  10p 10p 500p  1020p)

* setup the transient analysis
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot A0 A1 S X
.endc

.end
