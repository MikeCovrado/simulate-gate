
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulses for A0, A1 and S
*           pulse(V1  V2  TD    TR  TF  PW    PER)
Va0 A0 VGND pulse(0   1.8 1000p 10p 10p 1000p 2000p)
Va1 A1 VGND pulse(1.8 0   1000p 10p 10p 1000p 2000p)
Vs  S  VGND pulse(0   1.8  500p 10p 10p 2000p 4000p)

* setup the transient analysis
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot A0 A1
plot S
plot X
.endc

.end
